module and_gate (a,b,y);
	input a,b;
	output y;
	and g1(y,a,b);
endmodule

